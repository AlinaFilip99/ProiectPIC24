----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    13:50:48 03/17/2020 
-- Design Name: 
-- Module Name:    ROM32x32 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity ROM32x24 is
    Port ( Addr : in  STD_LOGIC_VECTOR (4 downto 0);
           Data : out  STD_LOGIC_VECTOR (23 downto 0));
end ROM32x24;

architecture Behavioral of ROM32x24 is
  type tROM is array (0 to 31) of STD_LOGIC_VECTOR (23 downto 0);
  
   constant ROM : tROM :=(
	             x"000001",-- 0000 0000 0000 0000 0000 0001
					 x"000002",-- 0000 0000 0000 0000 0000 0010
					 x"000004",-- 0000 0000 0000 0000 0000 0100
					 x"000008",-- 0000 0000 0000 0000 0000 1000
					 x"000010",-- 0000 0000 0000 0000 0001 0000
					 x"000020",-- 0000 0000 0000 0000 0010 0000
					 x"000040",-- 0000 0000 0000 0000 0100 0000
					 x"000080",-- 0000 0000 0000 0000 1000 0000
					 x"000100",-- 0000 0000 0000 0001 0000 0000
					 x"000200",-- 0000 0000 0000 0010 0000 0000
					 x"000400",-- 0000 0000 0000 0100 0000 0000
					 x"000800",-- 0000 0000 0000 1000 0000 0000
					 x"001000",-- 0000 0000 0001 0000 0000 0000
					 x"002000",-- 0000 0000 0010 0000 0000 0000
					 x"004000",-- 0000 0000 0100 0000 0000 0000
					 x"008000",-- 0000 0000 1000 0000 0000 0000
					 x"010000",-- 0000 0001 0000 0000 0000 0000
					 x"020000",-- 0000 0010 0000 0000 0000 0000
					 x"040000",-- 0000 0100 0000 0000 0000 0000
					 x"080000",-- 0000 1000 0000 0000 0000 0000
					 x"100000",-- 0001 0000 0000 0000 0000 0000
					 x"200000",-- 0010 0000 0000 0000 0000 0000
					 x"400000",-- 0100 0000 0000 0000 0000 0000
					 x"800000",-- 1000 0000 0000 0000 0000 0000
					 x"000000",-- 0000 0000 0000 0000 0000 0000
					 x"000000",-- 0000 0000 0000 0000 0000 0000
					 x"000000",-- 0000 0000 0000 0000 0000 0000
					 x"000000",-- 0000 0000 0000 0000 0000 0000
					 x"000000",-- 0000 0000 0000 0000 0000 0000
					 x"000000",-- 0000 0000 0000 0000 0000 0000
					 x"000000",-- 0000 0000 0000 0000 0000 0000
					 x"000000" );-- 0000 0000 0000 0000 0000 0000
					 
begin

    Data <= ROM(conv_integer(Addr));--Addr este PC(7:3)

end Behavioral;

